entity multiplexer is
port (
    i0, i1, i2, i3, a0, a1: in std_logic;
    x: out std_logic
);
end multiplexer;

architecture arq of multiplexer is
begin
    -- código aqui
end multiplexer
